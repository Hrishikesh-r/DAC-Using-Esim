* C:\Users\91990\AppData\Roaming\SPB_Data\eSim-Workspace\Switch_A\Switch_8A.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 09/30/21 11:38:56
.lib "sky130_fd_pr/models/sky130.lib.spice" tt

* Sheet Name: /
xM1  Vdd digital_Input Net-_M1-Pad3_ Vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5		
xM5  Net-_M1-Pad3_ digital_Input GND GND sky130_fd_pr__nfet_01v8 w=.42 l=.5		
xM2  Vdd Net-_M1-Pad3_ Net-_M2-Pad3_  Vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5		
xM6  Net-_M2-Pad3_ Net-_M1-Pad3_ GND GND sky130_fd_pr__nfet_01v8 w=.42 l=.5		
xM3   Vin_1 Net-_M1-Pad3_ Vout  Vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5		
xM7   Vout Net-_M1-Pad3_  Vin_2 GND sky130_fd_pr__nfet_01v8 w=.42 l=.5		
xM4   Vout Net-_M2-Pad3_  Vin_1 GND sky130_fd_pr__nfet_01v8 w=.42 l=.5		
xM8   Vin_2 Net-_M2-Pad3_  Vout  Vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5		

Vdd Vdd 0 3.3
Vin_1 Vin_1  0 2.5
Vin_2 Vin_2 0 2
Vd0 digital_Input 0 pulse(0 1.8 0s 0s 0s 5us 10us) 


.tran 0.1us 40us

.control
run

plot V(Vin_1) V(Vin_2) V(digital_Input) v(Vout) 


.endc

.end
